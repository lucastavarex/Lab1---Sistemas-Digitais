-------------- DATA: 22/06/2022                        --------------
-------------- AUTOR: LUCAS TAVARES DA SILVA FERREIRA  --------------
-------------- DRE: 120152739                          --------------
-------------- TÍTULO: TRABALHO 1 DE LABORATÓRIO       --------------
-------------- DISCIPLINA: SISTEMAS DIGITAIS           --------------
-------------- PROFESSOR: ROBERTO PACHECO              --------------


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADOR4 IS 
    PORT( 
		A, B: IN STD_LOGIC_VECTOR (3 DOWNTO 0);  -- VETORES DE ENTRADA DE 4 BITS A SEREM SOMADOS
		CARRY_IN: IN STD_LOGIC;                  -- CARRY
		SOMA: OUT STD_LOGIC_VECTOR (3 DOWNTO 0); -- RESULTADO
		CARRY_OUT,OVERFLOW: OUT STD_LOGIC        -- FLAGS DO RESULTADO 
		
            );
END SOMADOR4;

ARCHITECTURE DADOS OF SOMADOR4 IS
SIGNAL COUT,S,SOMA1,SOMA2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL X1, X2, X3, X4,X5,X6,X7,X8 : STD_LOGIC;


COMPONENT SOMADOR IS -- SOMADOR PARA CADA BIT
PORT ( 
A, B, CARRY_IN : IN STD_LOGIC;
SOMA, CARRY_OUT: OUT STD_LOGIC
);
END COMPONENT SOMADOR;



    BEGIN
        -- LÓGICA DE COMO FUNCIONA A SOMA 
        ADD0: SOMADOR PORT MAP(A(0), B(0), CARRY_IN, SOMA1(0), COUT(0));
        ADD1: SOMADOR PORT MAP(A(1), B(1), COUT(0), SOMA1(1), COUT(1)); -- CIN É O COUT DA OP ANTERIOR
        ADD2: SOMADOR PORT MAP(A(2), B(2), COUT(1), SOMA1(2), COUT(2));
        ADD3: SOMADOR PORT MAP(A(3), B(3), COUT(2), SOMA1(3), COUT(3));
     
    -- COMO OS NUMEROS A SEREM SOMADOS ESTÃO NO SISTEMA
    -- DE COMPLEMENTO DE 2 , TEREMOS QUE TRATÁ-LOS!

    X1 <= A(3) XNOR B(3);                          -- CASO TENHAM SINAIS IGUAIS
    X2 <= A(3) XOR B(3);                           -- CASO TENHAM SINAIS DIFERENTES
    X3 <= A(3) AND B(3);                           -- CASO AMBOS SEJAM NEGATIVOS
    X4 <= (NOT A(3)) AND (NOT B(3));               -- CASO AMBOS SEJAM POSITIVOS
    SOMA(3) <= (X1 AND A(3)) OR (X2 AND SOMA1(3)); -- FLAG DE SINAL SAI CERTO MESMO SE TIVER OVERFLOW
    SOMA(2) <= SOMA1(2);
	 SOMA(1) <= SOMA1(1);
	 SOMA(0) <= SOMA1(0);
    CARRY_OUT <=( X1 AND COUT(2)); -- SÓ TEM COUT SE OS SINAIS FOREM IGUAIS
    OVERFLOW <= (COUT(2) AND X4) OR (X3 AND (NOT(COUT(2)))); -- PARA O OVERFLOW, VAI DEPENDER SE OS SINAIS SÃO IGUAIS E 
                                                             -- SE ESTAMOS SOMANDO NÚMEROS NEGATIVOS OU POSITIVOS.
   
END DADOS;
