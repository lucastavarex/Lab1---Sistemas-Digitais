-------------- DATA: 22/06/2022                        --------------
-------------- AUTOR: LUCAS TAVARES DA SILVA FERREIRA  --------------
-------------- DRE: 120152739                          --------------
-------------- TÍTULO: TRABALHO 1 DE LABORATÓRIO       --------------
-------------- DISCIPLINA: SISTEMAS DIGITAIS           --------------
-------------- PROFESSOR: ROBERTO PACHECO              --------------


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUBTRADOR4 IS 
    PORT( 
		NA, NB: IN STD_LOGIC_VECTOR (3 DOWNTO 0) ;
		S: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0) ;
		SUBT: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		CARRY_OUT,OVERFLOW: OUT STD_LOGIC
            );
END SUBTRADOR4;

ARCHITECTURE DADOS OF SUBTRADOR4 IS
SIGNAL PSUB,X,Y : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
CONSTANT CC : STD_LOGIC :='1';  --  CIN = 1 PARA O COMPLEMENTO DE 2
SIGNAL COUT,OVRF : STD_LOGIC;



COMPONENT SOMADOR4 IS
PORT ( 
A, B: IN STD_LOGIC_VECTOR (3 DOWNTO 0); 
CARRY_IN: IN STD_LOGIC;
SOMA: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
CARRY_OUT,OVERFLOW: OUT STD_LOGIC
);
END COMPONENT SOMADOR4;

BEGIN
 
S <= NOT NB; -- RECEBE B BARRADO PARA O COMPLEMENTO DE 2

ADD : SOMADOR4 PORT MAP (NA, S, CC,SUBT,CARRY_OUT,OVERFLOW); -- FAZ A SOMA EM C2 ENTRE A E B NEGADO.
	 

END DADOS;